class MemScoreboard;

endclass
class AxiLiteDriver;
    
endclass
package axi_lite_sim;
    `include "./include/memory_transaction.sv"
    `include "./include/mem_active_driver.sv"
    `include "./include/mem_reactive_driver.sv"
endpackage

`timescale 1ns/1ps

class control;
    bit running;
endclass //control